
.param    P1_POS   = 0.9   ;Sweep
.param    P2_POS   = 0.9   ;Distortion
.param    MODE   = 1        ;Clip mode
.param    P3_POS   = 1   ;Filter
.param    P4_POS   = 0.9   ;Output volume

****************  GLOBAL SOURCES  ******************************************
VCC       VCC      0            DC 9
VIN       IN       0            SIN(0 50m 500)

****************  VIRTUAL HALF‑SUPPLY  *************************************
R10       VCC      VB           100k
R11       VB       0            100k
C13       VB       0            47u
C11       VCC      0            100u
C12       VCC      0            100n

****************  INPUT / PRE‑FILTER  **************************************
RPD       IN       0            2.2Meg
C1        IN       NIN          22n
R1        NIN      VB           1Meg
R2        NIN      AP1_Y        1k
C2        AP1_Y    0            1n

****************  SWEEP  (P1 – 1 kB)  **************************************
*.param    P1_POS   = 0.50
R3        AN1_Y    P1_A         47
RP1_A     P1_A     P1_W         {1k * P1_POS}
RP1_B     P1_W     P1_B         {1k * (1-P1_POS)}
RSHORT_P1 P1_B     P1_W         1u
C5        P1_B     0            2.2u

****************  OP‑AMP GAIN NETWORK  *************************************
R4        AN1_Y    NRKM1            560
C6        NRKM1    0            4.7u
*.param    P2_POS   = 0.50
*RP2_A     AN1_Y    P2_W         {100k * P2_POS}
*RP2_B     P2_W     AO1_Y        {100k * (1-P2_POS)}
RP2_A     AN1_Y    AO1_Y         {100k * P2_POS}
C4        AN1_Y    AO1_Y        100p
*XU1       AP1_Y    AN1_Y        AO1_Y      OP07      ;library subckt
XU1       AP1_Y    AN1_Y    VCC   0    AO1_Y      OP07      ;library subckt

****************  CLIPPING & MODE SWITCH  **********************************
C7        AO1_Y    CLIP_IN      4.7u
C14       AO1_Y    CLIP_IN      1u
R5        CLIP_IN  CLIP_SW      1k

*.param    MODE   = 1
BVCTL1    VCTL1    0            V={MODE}
BVCTL2    VCTL2    0            V={1-MODE}
S_MODE1   CLIP_SW  CLIP_CENT    VCTL1 0 SWMOD
S_MODE2   CLIP_SW  CLIP_PAIR    VCTL2 0 SWMOD

*diode arrays
D2        CLIP_PAIR 0           D1N914
D3        0         CLIP_PAIR   D1N914
D4        CLIP_CENT N_D4D5      D1N914
D5        N_D4D5    0           D1N914
D6        CLIP_CENT N_D6D7      D1N914
D7        N_D6D7    0           D1N914
D8        CLIP_CENT 0           D1N914   ;LED pair substituted with Si
D9        0         CLIP_CENT   D1N914
*rkmoore checked to here.  
****************  FILTER  (P3 – 100 kA)  ***********************************
*.param    P3_POS   = 0.50

*rkmoore: Is this next section hard-coded to the second switch position?
*left lug (P3_A) is CLIP_CENT, right lug (P3_B) feeds R6; wiper is P3_W.
RP3_A     CLIP_CENT P3_W        {100k * P3_POS}
RP3_B     P3_W      P3_B        {100k * (1-P3_POS)}
RSHORT_P3 CLIP_CENT P3_W        1u              ;lug‑3 ↔ wiper short as per PCB

R6        P3_B     BUF_IN       1.5k
C8        BUF_IN   0            3.3n
C9        BUF_IN   G1           22n
*R7        BUF_IN   0            1Meg
R7        G1       0            1Meg

****************  J‑FET OUTPUT BUFFER  *************************************
*Q1        D1       G1       S1      J2N5457      ;D G S
J1        D1       G1       S1      J2N5457      ;D G S
RD1       D1       VCC          1u               ;wire Drain → VCC
R8        S1       0            10k
C10       S1       VOUT_IN      1u

****************  VOLUME  (P4 – 100 kA)  ***********************************
*.param    P4_POS   = 0.75
RP4_A     VOUT_IN  P4_W         {100k * P4_POS}
RP4_B     P4_W     0            {100k * (1-P4_POS)}
R_ALIAS   OUT      P4_W         1u               ;OUT node alias

****************  ANALYSES  ************************************************
*.op
*.tran     0 20m 0 10u
*.tran     2u 100m 80m


****************  MODELS  (alphabetical)  **********************************
.model    D1N914  D
.model    J2N5457 NJF(Beta=1.72m Vto=-2.03 Lambda=50m Rs=1 Rd=1)
.model    SWMOD   SW(Ron=0.1 Roff=1e9 Vt=0.5 Vh=0.1)
.subckt IDEALOPAMP 1 2 6         ; +, –, out
EGAIN  7 0  1 2 1e6
Rout   6 7  10
Cout   7 0  1p
.ends  IDEALOPAMP

****************  LIBRARIES  ***********************************************
*.include  OP07.cir          *adjust path to ngspice/examples if needed

* 
* Linear Technology OP07 op amp model
* Written: 08-24-1989 12:35:59 Type: Bipolar npn input, internal comp.
* Typical specs: 
* Vos=3.0E-05, Ib=1.0E-09, Ios=4.0E-10, GBP=6.0E+05Hz, Phase mar.= 70 deg, 
* SR(+)=2.5E-01V/us, SR(-)=2.4E-01V/us, Av= 114 dB, CMMR= 126 dB, 
* Vsat(+)=2.00V, Vsat(-)=2.00V, Isc=+/-25.0mA, Iq=2500uA
* (input differential mode clamp active)
* 
* Connections: + - V+V-O 
.subckt OP07 3 2 7 4 6
* input
rc1 7  80 8.842E+03
rc2 7  90 8.842E+03
q1  80 102 10 qm1 
q2  90 103 11 qm2 
rb1  2   102 5.000E+02
rb2  3   103 5.000E+02
ddm1 102 104 dm2 
ddm3 104 103 dm2 
ddm2 103 105 dm2 
ddm4 105 102 dm2 
c1  80 90 5.460E-12
re1 10 12 1.948E+03
re2 11 12 1.948E+03
iee 12 4  7.502E-06
re  12 0  2.666E+07
ce  12 0  1.579E-12
* intermediate 
gcm 0  8  12 0  5.668E-11
ga  8  0  80 90 1.131E-04
r2  8  0  1.000E+05
c2  1  8  3.000E-11
gb  1  0  8  0  1.294E+03
* output 
ro1 1  6  2.575E+01
ro2 1  0  3.425E+01
rc  17 0  6.634E-06
gc  0  17 6  0  1.507E+05
d1  1  17 dm1 
d2  17 1  dm1 
d3  6  13 dm2 
d4  14 6  dm2 
vc  7  13 2.803E+00
ve  14 4  2.803E+00
ip  7  4  2.492E-03
dsub 4  7  dm2 
* models 
.model qm1 npn (is=8.000E-16 bf=3.125E+03)
.model qm2 npn (is=8.009E-16 bf=4.688E+03)
.model dm1 d   (is=1.486E-08)
.model dm2 d   (is=8.000E-16)
.ends OP07
* 
* - - - - - * fini OP07 * - - - - - * [oamm vn1 8/89]
**
*         (C) COPYRIGHT LINEAR TECHNOLOGY CORPORATION 1990
*                       All rights reserved.
* 
*   Linear Technology Corporation hereby grants the users of this
* macromodel a non-exclusive, nontransferrable license to use this
*            macromodel under the following conditions:
* 
* The user agrees that this macromodel is licensed from Linear
* Technology and agrees that the macromodel may be used, loaned,
* given away or included in other model libraries as long as this
* notice and the model in its entirety and unchanged is included.
* No right to make derivative works or modifications to the
* macromodel is granted hereby.  All such rights are reserved.
* 
* This model is provided as is.  Linear Technology makes no
* warranty, either expressed or implied about the suitability or
* fitness of this model for any particular purpose.  In no event
* will Linear Technology be liable for special, collateral,
* incidental or consequential damages in connection with or arising
* out of the use of this macromodel.  It should be remembered that
* models are a simplification of the actual circuit.
* 
* Linear Technology reserves the right to change these macromodels
* without prior notice.  Contact Linear Technology at 1630 McCarthy
* Blvd., Milpitas, CA, 95035-7487 or telephone 408/432-1900 for
* datasheets on the actual amplifiers or the latest macromodels.
* 
* ----------------------------------------------------------------------- *
**.tran 2u 100m 80m
**.op
**.control
**  run
**  plot v(IN) v(OUT)
**.endc
**.end

.tran 2u 100m 80m
.op
.control
  run
  *plot v(IN) v(OUT)
 ** plot v(OUT)
 * plot db(OUT)
 print OUT
 quit
.endc
.end
