*ProcoRatV0.cir
*------------------------------------------------------------
* Pro Co RAT distortion (Aion Helios) – ngspice netlist
* 9 V single-rail; rail-protection / conditioning removed
*------------------------------------------------------------

*--- GLOBAL SOURCES ---
VCC   VCC   0              DC 9
VIN   IN    0              SIN(0 50m 500)

*--- REFERENCE (VB ≈ 4.5 V) ---
R10   VCC   VB             100k
R11   VB    0              100k
C13   VB    0              47u      ;virtual-ground filter
C11   VCC    0              100u
C12   VCC    0              100n

*--- INPUT / PRE-FILTER ---
RPD   IN    0              2.2Meg
C1    IN    NIN_P          22n
R2    NIN_P VB             1Meg
R3    NIN_P AN1_Y          1k
C2    AN1_Y 0              1n

*--- OP-AMP (ideal vcvs, OP07 comp cap omitted) ---
EOP   AO1_Y 0   AN1_Y AP1_Y  1e6
AP1_Y VB                   ;non-inverting input is VB

*--- FEEDBACK / GAIN (DIST pot) ---
R4    AN1_Y NF             47
R5    AN1_Y NF             560
C5    NF    0              2.2u
C6    NF    0              4.7u
C4    NF    AO1_Y          100p

.param DIST_POS=0.5        ;0=minimum gain, 1=max
P_DIST_A NF  P_DIST_W      {100k*DIST_POS}
P_DIST_B P_DIST_W AO1_Y    {100k*(1-DIST_POS)}

*--- CLIPPING STAGE ---
C7    AO1_Y NCLIP_IN       4.7u
R6    NCLIP_IN NCLIP       1k
D2    NCLIP   0            D1N914
D3    0       NCLIP        D1N914

*--- TONE (FILTER pot wired “reversed” as in RAT) ---
.param FILTER_POS=0.5
P_FIL_A NCLIP N_FIL_W      {100k*FILTER_POS}
P_FIL_B N_FIL_W NCLIP      {100k*(1-FILTER_POS)}
R7     N_FIL_W NOUT_BUF_G  1.5k
C8     NOUT_BUF_G 0        3.3n

*--- OUTPUT BUFFER (2N5485 source follower) ---
C9    NOUT_BUF_G G1        22n
R8    G1     0             1Meg
Q1    D1     G1  S1        J2N5485
D1    VCC                  ;drain at 9 V
R9    S1     0             10k
C10   S1     N_VOL_IN      1u

*--- VOLUME pot ---
.param VOL_POS=0.75        ;0=mute, 1=max
P_VOL_A N_VOL_IN  VOUT     {100k*VOL_POS}
P_VOL_B VOUT      0        {100k*(1-VOL_POS)}

*--- ANALYSES ---
.op
.tran 0 20m 0 10u

*--- MODELS (alphabetical) ---
.model D1N914 D
.model J2N5485 NJF(VTO=-2 BETA=3.5m LAMBDA=10m)
.control
  * quick sanity check
  * 100 mVp 1 kHz sine
  *vin IN 0 SIN(0 0.1 1k)

  * comment the next two lines and uncomment the .ac if you’d rather sweep
  *tran 5u 100m
  tran 2u 100m 80m
  plot v(IN) v(OUT)

  *ac dec 30 20 20k
.endc
.end
