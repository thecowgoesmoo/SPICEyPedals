
.param    P1_POS   = 0.98   ;Drive
.param    P2_POS   = 0.98   ;Tone
.param    P3_POS   = 0.98   ;Level

*IbanezTS9.cir
*-------------------------------------------------------------
*  Stratus / Ibanez TS-9 audio core – NGSPICE .cir
*  Default stimulus : 500 Hz, 50 mVpk sine
*  Transient plot   : 80 ms → 100 ms, 2 µs step
*-------------------------------------------------------------
* SIGNAL SOURCE ------------------------------------------------
vin  IN  0  SIN(0 0.05 500)      ; 50 mVpk, 500 Hz

* SUPPLY & VIRTUAL MID-RAIL -----------------------------------
VCC   9V  0   DC 9
R16   9V  VB  10k
R17   VB  0   10k
C11   VB  0   47u
C12   VB  0   100n
C10   9V  0   100u
C13   9V  0   100n

* INPUT NETWORK ------------------------------------------------
C1   IN  NN1  22n
RPD  IN  0   2.2Meg
R1   NN1 B1  1k
R2   B1  VB  510k                ; bias to mid-rail

*Buffer stage
Q1 9V B1 E1 2N5088
R3 E1 0 10k

* OP-AMP A  (DISTORTION) --------------------------------------
C2 E1 N1_1 1u
XU1A N1_1 N1_2 A1_1  IDEALOPAMP        ; non-inv, inv, out
R4 VB   N1_1 10k

C3 A1_1 N1_2 47p
D2 A1_1  N1_2  D1N914
D3 N1_2  A1_1  D1N914
***RD2 A1_1 N1_2  1k
***RD3 N1_2  A1_1 1k
**D4 A1_1 NN1 D1N914
**D5 NN1 N1_2 D1N914
**D7 NN2 A1_1 D1N914
**D6 N1_2 NN2 D1N914
D8 A1_1 N1_2  LED1
D9 N1_2 A1_1  LED1
***RD8 A1_1 N1_2  1k
***RD9 N1_2 A1_1  1k
C4 N1_2 NN6 47n
R5 NN6  VB  4.7k

*Drive pot in a middle position
*RDRV A1_1 N1_2 300k
RDRV A1_1 N1_2 {P1_POS*500k+50k} 

*rkmoore checked to here  

* Drive pot (500 kΩ) centred → two 250 kΩ sections

* Symmetrical Si clipping diodes (stock position)

* COUPLING TO TONE STACK --------------------------------------
R7 A1_1 N2_1 1k
R8 N2_1 VB   10k
C5 N2_1 0    220n
C6 NT   NN5  220n                ; mid-hump 
R9 NN5  0    220

* TONE POT (20 kΩ W pot, centre)
*RT_T NT  N2_2   10k
*RT_B N2_1  NT   10k                 ; wiper node = NT
RT_T NT  N2_2   {(1-P2_POS)*10k}
RT_B N2_1  NT   {P2_POS*10k}                 ; wiper node = NT
*rkmoore double check to here
* OP-AMP B  (BUFFER / LEVEL) ----------------------------------
* Unity-gain non-inverting buffer biased at VB
XU1B N2_1  N2_2  A2_1  IDEALOPAMP
R10 A2_1 N2_2 1k
C7  A2_1 NN3 1u
R11 NN3 VOL_TOP 1k

* LEVEL POT (100 kΩ A pot, centre)
*RV_T VOL_TOP VOL_W 1k
*RV_B VOL_W   VB    99k
RV_T VOL_TOP VOL_W {(1-P3_POS)*10k}
RV_B VOL_W   VB    {P3_POS*10k}

*Output buffer
C8  VOL_W B2  100n
R12 B2    VB  510k
Q2  9V    B2  E2 2N5088
R13 E2    0   10k
R14 E2    NN4 100
C9  NN4   OUT 1u
R15 OUT   0   10k

*-------------------------------------------------------------
* DEVICE MODELS ------------------------------------------------
*.model D1N914 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n Iave=200m Vpk=75)
.model 2N5088 NPN (BF=300 IS=5e-15 VAF=100)
.model D1N914 D(IS=2.52e-9 RS=10 CJO=2pF N=1.7 BV=100)
.MODEL LED1 D (
+ IS=93.2P  N=1.78 BV=4  IBV=10U RS=0.15  VJ=0.7  
+ LED  IF=40m  trr=3u )
* Simple wide-band ideal op-amp (good enough for time-domain)
.subckt IDEALOPAMP 1 2 6         ; +, –, out
EGAIN  7 0  1 2 1e6
Rout   6 7  10
Cout   7 0  1p
.ends  IDEALOPAMP

*-------------------------------------------------------------
* ANALYSIS -----------------------------------------------------
*.tran 2u 100m 80m
*.op
*.control
*  run
*  plot v(IN) v(OUT)
*.endc
*.end

.tran 2u 100m 80m
.op
.control
  run
  *plot v(IN) v(OUT)
 ** plot v(OUT)
 * plot db(OUT)
 print OUT
 quit
.endc
.end
