
.param    P1_POS   = 0.98   ;Harmonics
.param    P2_POS   = 0.99   ;Balance

*---------------------------------------------------------------------------
*  AION “PARTICLE”  –  Interfax Harmonic Percolator (ALBINI spec, 9 V)
*---------------------------------------------------------------------------

***** SUPPLY & POWER FILTER ***********************************************
VRAW    9VRAW     0           DC 9             ; battery / adaptor
vin     IN        0           SIN(0 0.05 500)

***** INPUT / “HARMONICS” POT *********************************************
* 100 k log pot wired as variable series resistor, full-up by default

*RP2_A     AN1_Y    P2_W         {100k * P2_POS}
*RP2_B     P2_W     AO1_Y        {100k * (1-P2_POS)}

*RHPOT_T IN      HARM_W     1
*RHPOT_B HARM_W  0          99k               ; 1 Ω + 99 k ≈ 100 kA @ max

RHPOT_T IN      HARM_W     {100k * (1-P1_POS)}
RHPOT_B HARM_W  0          {100k * P1_POS}               

* 47 n coupling cap into PNP base
C2      HARM_W  B_PNP      47n

***** BIAS & FEEDBACK NETWORK *********************************************
R1      B_PNP    C_PNP      51k                ; Albini input bias to GND
R3      C_NPN    B_NPN      3.9Meg             ; positive feedback
R4      9VRAW     C_NPN     91k                ; Q1 base-to-collector bias

***** TRANSISTOR PAIR *****************************************************
* Node legend:  C  B  E   (arrow is on emitter – both emitters share node J)
Q1      C_PNP   B_PNP   J          2N404A_PNP
Q2      C_NPN   B_NPN   J          2N3904_NPN

* Collector loads
R2      C_PNP     0     91k                  ; Albini value
R5      BAL_TOP   D2AN  4.7k                 ; to ground per Albini schematic

* Shared emitter node bypass
C3      J        0          47u
C4      B_NPN    C_PNP     2.2u
***** SMALL SHAPING CAPS **************************************************
C1      HARM_W   0          100p                ; RF roll-off
C5      C_PNP    0          1.5n                ; mid-boost contour

***** CLIPPING SECTION – “MODE” SWITCH ************************************
*     SPDT centre-off wired as three positions:
*     - Ge pair (D2,D3)    - Si pair (D4–D7 in series pairs)   - None
D2      D2AN     0          D_GE
D3      0        BAL_TOP    D_GE
*D4      BAL_TOP  CLIP1      1N914
*D5      CLIP1    0          1N914
*D6      0        CLIP2      1N914
*D7      CLIP2    BAL_TOP    1N914
*SCLP_G  C_NPN   0      CLP_SW  VCTL_G         ; Ge position
*SCLP_S  C_NPN   0      CLP_SW  VCTL_S         ; Si position
* VCTL_G / VCTL_S are ideal logic sources that you toggle 1=>0 to pick the branch.
* For casual sims just comment one “S” device to select the diode set.

.model CLP_SW SW(Ron=0.01 Roff=1e9 Vt=0.5 Vh=0.1)  ; perfect-ish switch model

***** OUTPUT / “BALANCE” POT **********************************************
C6      C_NPN    BAL_TOP    100n               ; 100 nF output coupling
*RBAL_T  BAL_TOP  OUT        1
*RBAL_B  OUT      0          49.0k              ; 50 kA at full clockwise
RBAL_T  BAL_TOP  OUT        {50k * (1-P2_POS)}
RBAL_B  OUT      0          {50k * P2_POS}              ; 50 kA at full clockwise

***** DEVICE MODELS (quick generic) ***************************************
.model 2N404A_PNP PNP(BF=50  IS=1e-9  VAF=60)
.model 2N3904_NPN NPN(BF=180 IS=5e-15 VAF=100)
.model D_GE D(IS=5u RS=2 N=1.7 CJO=20p)
.model D1N5817 D(IS=35u N=1.1 RS=0.05 CJO=110p TT=10n)
.model 1N914 D (Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n Iave=200m Vpk=75)

*---------------------------------------------------------------------------
*.control
*  * Small-signal frequency sweep
*  *ac dec 30 20 20k
*  *plot vdb(IN) vdb(OUT)
*  * Transient test – 200 mVp, 500 Hz sine into full-CW Harmonics  
*  tran 2u 100m 80m
*  *plot v(IN) v(OUT)
*plot v(OUT)
**plot v(IN) vs v(OUT)
**plot v(OUT) vs v(IN)
*.endc
*.end

.tran 2u 100m 80m
.op
.control
  run
  *plot v(IN) v(OUT)
 ** plot v(OUT)
 * plot db(OUT)
 print OUT
 quit
.endc
.end


